// master_nios_multiple_slave.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module master_nios_multiple_slave (
		input  wire [31:0] aip_up_0_aip_dataout, //   aip_up_0.aip_dataout
		input  wire        aip_up_0_aip_int,     //           .aip_int
		output wire [4:0]  aip_up_0_aip_config,  //           .aip_config
		output wire [31:0] aip_up_0_aip_datain,  //           .aip_datain
		output wire        aip_up_0_aip_read,    //           .aip_read
		output wire        aip_up_0_aip_write,   //           .aip_write
		output wire        aip_up_0_core_int,    //           .core_int
		output wire        aip_up_0_aip_start,   //           .aip_start
		input  wire        clk_clk,              //        clk.clk
		input  wire [7:0]  int_ip_s0_export,     //  int_ip_s0.export
		output wire [9:0]  leds_export,          //       leds.export
		input  wire [31:0] port_s0_aip_dataout,  //    port_s0.aip_dataout
		input  wire        port_s0_aip_int,      //           .aip_int
		output wire [4:0]  port_s0_aip_config,   //           .aip_config
		output wire [31:0] port_s0_aip_datain,   //           .aip_datain
		output wire        port_s0_aip_read,     //           .aip_read
		output wire        port_s0_aip_write,    //           .aip_write
		output wire        port_s0_core_int,     //           .core_int
		output wire        port_s0_aip_start,    //           .aip_start
		input  wire [31:0] port_s1_aip_dataout,  //    port_s1.aip_dataout
		input  wire        port_s1_aip_int,      //           .aip_int
		output wire [4:0]  port_s1_aip_config,   //           .aip_config
		output wire [31:0] port_s1_aip_datain,   //           .aip_datain
		output wire        port_s1_aip_read,     //           .aip_read
		output wire        port_s1_aip_write,    //           .aip_write
		output wire        port_s1_core_int,     //           .core_int
		output wire        port_s1_aip_start,    //           .aip_start
		input  wire [31:0] port_s2_aip_dataout,  //    port_s2.aip_dataout
		input  wire        port_s2_aip_int,      //           .aip_int
		output wire [4:0]  port_s2_aip_config,   //           .aip_config
		output wire [31:0] port_s2_aip_datain,   //           .aip_datain
		output wire        port_s2_aip_read,     //           .aip_read
		output wire        port_s2_aip_write,    //           .aip_write
		output wire        port_s2_core_int,     //           .core_int
		output wire        port_s2_aip_start,    //           .aip_start
		input  wire        reset_reset_n,        //      reset.reset_n
		input  wire        spi_MISO,             //        spi.MISO
		output wire        spi_MOSI,             //           .MOSI
		output wire        spi_SCLK,             //           .SCLK
		output wire        spi_SS_n,             //           .SS_n
		input  wire        start_up_0_export,    // start_up_0.export
		input  wire        uart_rxd,             //       uart.rxd
		output wire        uart_txd              //           .txd
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [18:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [18:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_aip_up_0_avalon_slave_0_chipselect;        // mm_interconnect_0:aip_uP_0_avalon_slave_0_chipselect -> aip_uP_0:chipselect
	wire  [31:0] mm_interconnect_0_aip_up_0_avalon_slave_0_readdata;          // aip_uP_0:readdata -> mm_interconnect_0:aip_uP_0_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_aip_up_0_avalon_slave_0_address;           // mm_interconnect_0:aip_uP_0_avalon_slave_0_address -> aip_uP_0:address
	wire         mm_interconnect_0_aip_up_0_avalon_slave_0_read;              // mm_interconnect_0:aip_uP_0_avalon_slave_0_read -> aip_uP_0:read
	wire         mm_interconnect_0_aip_up_0_avalon_slave_0_write;             // mm_interconnect_0:aip_uP_0_avalon_slave_0_write -> aip_uP_0:write
	wire  [31:0] mm_interconnect_0_aip_up_0_avalon_slave_0_writedata;         // mm_interconnect_0:aip_uP_0_avalon_slave_0_writedata -> aip_uP_0:writedata
	wire         mm_interconnect_0_aip_1_avalon_slave_0_chipselect;           // mm_interconnect_0:aip_1_avalon_slave_0_chipselect -> aip_1:chipselect
	wire  [31:0] mm_interconnect_0_aip_1_avalon_slave_0_readdata;             // aip_1:readdata -> mm_interconnect_0:aip_1_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_aip_1_avalon_slave_0_address;              // mm_interconnect_0:aip_1_avalon_slave_0_address -> aip_1:address
	wire         mm_interconnect_0_aip_1_avalon_slave_0_read;                 // mm_interconnect_0:aip_1_avalon_slave_0_read -> aip_1:read
	wire         mm_interconnect_0_aip_1_avalon_slave_0_write;                // mm_interconnect_0:aip_1_avalon_slave_0_write -> aip_1:write
	wire  [31:0] mm_interconnect_0_aip_1_avalon_slave_0_writedata;            // mm_interconnect_0:aip_1_avalon_slave_0_writedata -> aip_1:writedata
	wire         mm_interconnect_0_aip_2_avalon_slave_0_chipselect;           // mm_interconnect_0:aip_2_avalon_slave_0_chipselect -> aip_2:chipselect
	wire  [31:0] mm_interconnect_0_aip_2_avalon_slave_0_readdata;             // aip_2:readdata -> mm_interconnect_0:aip_2_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_aip_2_avalon_slave_0_address;              // mm_interconnect_0:aip_2_avalon_slave_0_address -> aip_2:address
	wire         mm_interconnect_0_aip_2_avalon_slave_0_read;                 // mm_interconnect_0:aip_2_avalon_slave_0_read -> aip_2:read
	wire         mm_interconnect_0_aip_2_avalon_slave_0_write;                // mm_interconnect_0:aip_2_avalon_slave_0_write -> aip_2:write
	wire  [31:0] mm_interconnect_0_aip_2_avalon_slave_0_writedata;            // mm_interconnect_0:aip_2_avalon_slave_0_writedata -> aip_2:writedata
	wire         mm_interconnect_0_aip_0_avalon_slave_0_chipselect;           // mm_interconnect_0:aip_0_avalon_slave_0_chipselect -> aip_0:chipselect
	wire  [31:0] mm_interconnect_0_aip_0_avalon_slave_0_readdata;             // aip_0:readdata -> mm_interconnect_0:aip_0_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_aip_0_avalon_slave_0_address;              // mm_interconnect_0:aip_0_avalon_slave_0_address -> aip_0:address
	wire         mm_interconnect_0_aip_0_avalon_slave_0_read;                 // mm_interconnect_0:aip_0_avalon_slave_0_read -> aip_0:read
	wire         mm_interconnect_0_aip_0_avalon_slave_0_write;                // mm_interconnect_0:aip_0_avalon_slave_0_write -> aip_0:write
	wire  [31:0] mm_interconnect_0_aip_0_avalon_slave_0_writedata;            // mm_interconnect_0:aip_0_avalon_slave_0_writedata -> aip_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_start_up_s1_chipselect;                    // mm_interconnect_0:start_uP_s1_chipselect -> start_uP:chipselect
	wire  [31:0] mm_interconnect_0_start_up_s1_readdata;                      // start_uP:readdata -> mm_interconnect_0:start_uP_s1_readdata
	wire   [1:0] mm_interconnect_0_start_up_s1_address;                       // mm_interconnect_0:start_uP_s1_address -> start_uP:address
	wire         mm_interconnect_0_start_up_s1_write;                         // mm_interconnect_0:start_uP_s1_write -> start_uP:write_n
	wire  [31:0] mm_interconnect_0_start_up_s1_writedata;                     // mm_interconnect_0:start_uP_s1_writedata -> start_uP:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [3:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_int_ip_s0_s1_chipselect;                   // mm_interconnect_0:int_IP_s0_s1_chipselect -> int_IP_s0:chipselect
	wire  [31:0] mm_interconnect_0_int_ip_s0_s1_readdata;                     // int_IP_s0:readdata -> mm_interconnect_0:int_IP_s0_s1_readdata
	wire   [1:0] mm_interconnect_0_int_ip_s0_s1_address;                      // mm_interconnect_0:int_IP_s0_s1_address -> int_IP_s0:address
	wire         mm_interconnect_0_int_ip_s0_s1_write;                        // mm_interconnect_0:int_IP_s0_s1_write -> int_IP_s0:write_n
	wire  [31:0] mm_interconnect_0_int_ip_s0_s1_writedata;                    // mm_interconnect_0:int_IP_s0_s1_writedata -> int_IP_s0:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                        // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                          // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                           // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                             // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                         // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                      // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                        // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                         // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                            // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                   // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                           // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                       // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         mm_interconnect_0_mem_data_s1_chipselect;                    // mm_interconnect_0:mem_data_s1_chipselect -> mem_data:chipselect
	wire  [31:0] mm_interconnect_0_mem_data_s1_readdata;                      // mem_data:readdata -> mm_interconnect_0:mem_data_s1_readdata
	wire  [11:0] mm_interconnect_0_mem_data_s1_address;                       // mm_interconnect_0:mem_data_s1_address -> mem_data:address
	wire   [3:0] mm_interconnect_0_mem_data_s1_byteenable;                    // mm_interconnect_0:mem_data_s1_byteenable -> mem_data:byteenable
	wire         mm_interconnect_0_mem_data_s1_write;                         // mm_interconnect_0:mem_data_s1_write -> mem_data:write
	wire  [31:0] mm_interconnect_0_mem_data_s1_writedata;                     // mm_interconnect_0:mem_data_s1_writedata -> mem_data:writedata
	wire         mm_interconnect_0_mem_data_s1_clken;                         // mm_interconnect_0:mem_data_s1_clken -> mem_data:clken
	wire         mm_interconnect_0_spi_0_spi_control_port_chipselect;         // mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_readdata;           // spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_0_spi_control_port_address;            // mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire         mm_interconnect_0_spi_0_spi_control_port_read;               // mm_interconnect_0:spi_0_spi_control_port_read -> spi_0:read_n
	wire         mm_interconnect_0_spi_0_spi_control_port_write;              // mm_interconnect_0:spi_0_spi_control_port_write -> spi_0:write_n
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_writedata;          // mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire         mm_interconnect_0_mem_program_s1_chipselect;                 // mm_interconnect_0:mem_program_s1_chipselect -> mem_program:chipselect
	wire  [31:0] mm_interconnect_0_mem_program_s1_readdata;                   // mem_program:readdata -> mm_interconnect_0:mem_program_s1_readdata
	wire  [15:0] mm_interconnect_0_mem_program_s1_address;                    // mm_interconnect_0:mem_program_s1_address -> mem_program:address
	wire   [3:0] mm_interconnect_0_mem_program_s1_byteenable;                 // mm_interconnect_0:mem_program_s1_byteenable -> mem_program:byteenable
	wire         mm_interconnect_0_mem_program_s1_write;                      // mm_interconnect_0:mem_program_s1_write -> mem_program:write
	wire  [31:0] mm_interconnect_0_mem_program_s1_writedata;                  // mm_interconnect_0:mem_program_s1_writedata -> mem_program:writedata
	wire         mm_interconnect_0_mem_program_s1_clken;                      // mm_interconnect_0:mem_program_s1_clken -> mem_program:clken
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // start_uP:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // int_IP_s0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // uart_0:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                    // spi_0:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [aip_0:resetn, aip_1:resetn, aip_2:resetn, aip_uP_0:resetn, irq_mapper:reset, leds:reset_n, mem_program:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset, start_uP:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [int_IP_s0:reset_n, jtag_uart_0:rst_n, mem_data:reset, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_translator_001:in_reset, spi_0:reset_n, timer_0:reset_n, uart_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [mem_data:reset_req, rst_translator_001:reset_req_in]

	avalon_aip_avalon_interface aip_0 (
		.address              (mm_interconnect_0_aip_0_avalon_slave_0_address),    //        avalon_slave_0.address
		.chipselect           (mm_interconnect_0_aip_0_avalon_slave_0_chipselect), //                      .chipselect
		.write                (mm_interconnect_0_aip_0_avalon_slave_0_write),      //                      .write
		.writedata            (mm_interconnect_0_aip_0_avalon_slave_0_writedata),  //                      .writedata
		.read                 (mm_interconnect_0_aip_0_avalon_slave_0_read),       //                      .read
		.readdata             (mm_interconnect_0_aip_0_avalon_slave_0_readdata),   //                      .readdata
		.resetn               (~rst_controller_reset_out_reset),                   //                 reset.reset_n
		.clk                  (clk_clk),                                           //                   clk.clk
		.i_aip_dataOut_export (port_s0_aip_dataout),                               // external_connection_1.aip_dataout
		.i_aip_int_export     (port_s0_aip_int),                                   //                      .aip_int
		.o_aip_config_export  (port_s0_aip_config),                                //                      .aip_config
		.o_aip_dataIn_export  (port_s0_aip_datain),                                //                      .aip_datain
		.o_aip_read_export    (port_s0_aip_read),                                  //                      .aip_read
		.o_aip_write_export   (port_s0_aip_write),                                 //                      .aip_write
		.o_core_int_export    (port_s0_core_int),                                  //                      .core_int
		.o_aip_start_export   (port_s0_aip_start)                                  //                      .aip_start
	);

	avalon_aip_avalon_interface aip_1 (
		.address              (mm_interconnect_0_aip_1_avalon_slave_0_address),    //        avalon_slave_0.address
		.chipselect           (mm_interconnect_0_aip_1_avalon_slave_0_chipselect), //                      .chipselect
		.write                (mm_interconnect_0_aip_1_avalon_slave_0_write),      //                      .write
		.writedata            (mm_interconnect_0_aip_1_avalon_slave_0_writedata),  //                      .writedata
		.read                 (mm_interconnect_0_aip_1_avalon_slave_0_read),       //                      .read
		.readdata             (mm_interconnect_0_aip_1_avalon_slave_0_readdata),   //                      .readdata
		.resetn               (~rst_controller_reset_out_reset),                   //                 reset.reset_n
		.clk                  (clk_clk),                                           //                   clk.clk
		.i_aip_dataOut_export (port_s1_aip_dataout),                               // external_connection_1.aip_dataout
		.i_aip_int_export     (port_s1_aip_int),                                   //                      .aip_int
		.o_aip_config_export  (port_s1_aip_config),                                //                      .aip_config
		.o_aip_dataIn_export  (port_s1_aip_datain),                                //                      .aip_datain
		.o_aip_read_export    (port_s1_aip_read),                                  //                      .aip_read
		.o_aip_write_export   (port_s1_aip_write),                                 //                      .aip_write
		.o_core_int_export    (port_s1_core_int),                                  //                      .core_int
		.o_aip_start_export   (port_s1_aip_start)                                  //                      .aip_start
	);

	avalon_aip_avalon_interface aip_2 (
		.address              (mm_interconnect_0_aip_2_avalon_slave_0_address),    //        avalon_slave_0.address
		.chipselect           (mm_interconnect_0_aip_2_avalon_slave_0_chipselect), //                      .chipselect
		.write                (mm_interconnect_0_aip_2_avalon_slave_0_write),      //                      .write
		.writedata            (mm_interconnect_0_aip_2_avalon_slave_0_writedata),  //                      .writedata
		.read                 (mm_interconnect_0_aip_2_avalon_slave_0_read),       //                      .read
		.readdata             (mm_interconnect_0_aip_2_avalon_slave_0_readdata),   //                      .readdata
		.resetn               (~rst_controller_reset_out_reset),                   //                 reset.reset_n
		.clk                  (clk_clk),                                           //                   clk.clk
		.i_aip_dataOut_export (port_s2_aip_dataout),                               // external_connection_1.aip_dataout
		.i_aip_int_export     (port_s2_aip_int),                                   //                      .aip_int
		.o_aip_config_export  (port_s2_aip_config),                                //                      .aip_config
		.o_aip_dataIn_export  (port_s2_aip_datain),                                //                      .aip_datain
		.o_aip_read_export    (port_s2_aip_read),                                  //                      .aip_read
		.o_aip_write_export   (port_s2_aip_write),                                 //                      .aip_write
		.o_core_int_export    (port_s2_core_int),                                  //                      .core_int
		.o_aip_start_export   (port_s2_aip_start)                                  //                      .aip_start
	);

	avalon_aip_avalon_interface aip_up_0 (
		.address              (mm_interconnect_0_aip_up_0_avalon_slave_0_address),    //        avalon_slave_0.address
		.chipselect           (mm_interconnect_0_aip_up_0_avalon_slave_0_chipselect), //                      .chipselect
		.write                (mm_interconnect_0_aip_up_0_avalon_slave_0_write),      //                      .write
		.writedata            (mm_interconnect_0_aip_up_0_avalon_slave_0_writedata),  //                      .writedata
		.read                 (mm_interconnect_0_aip_up_0_avalon_slave_0_read),       //                      .read
		.readdata             (mm_interconnect_0_aip_up_0_avalon_slave_0_readdata),   //                      .readdata
		.resetn               (~rst_controller_reset_out_reset),                      //                 reset.reset_n
		.clk                  (clk_clk),                                              //                   clk.clk
		.i_aip_dataOut_export (aip_up_0_aip_dataout),                                 // external_connection_1.aip_dataout
		.i_aip_int_export     (aip_up_0_aip_int),                                     //                      .aip_int
		.o_aip_config_export  (aip_up_0_aip_config),                                  //                      .aip_config
		.o_aip_dataIn_export  (aip_up_0_aip_datain),                                  //                      .aip_datain
		.o_aip_read_export    (aip_up_0_aip_read),                                    //                      .aip_read
		.o_aip_write_export   (aip_up_0_aip_write),                                   //                      .aip_write
		.o_core_int_export    (aip_up_0_core_int),                                    //                      .core_int
		.o_aip_start_export   (aip_up_0_aip_start)                                    //                      .aip_start
	);

	master_nios_multiple_slave_int_IP_s0 int_ip_s0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_int_ip_s0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_int_ip_s0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_int_ip_s0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_int_ip_s0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_int_ip_s0_s1_readdata),   //                    .readdata
		.in_port    (int_ip_s0_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                   //                 irq.irq
	);

	master_nios_multiple_slave_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	master_nios_multiple_slave_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	master_nios_multiple_slave_mem_data mem_data (
		.clk        (clk_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_mem_data_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_mem_data_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_mem_data_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_mem_data_s1_write),      //       .write
		.readdata   (mm_interconnect_0_mem_data_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_mem_data_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_mem_data_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                      // (terminated)
	);

	master_nios_multiple_slave_mem_program mem_program (
		.clk        (clk_clk),                                     //   clk1.clk
		.address    (mm_interconnect_0_mem_program_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_mem_program_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_mem_program_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_mem_program_s1_write),      //       .write
		.readdata   (mm_interconnect_0_mem_program_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_mem_program_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_mem_program_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req  (1'b0),                                        // (terminated)
		.freeze     (1'b0)                                         // (terminated)
	);

	master_nios_multiple_slave_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	master_nios_multiple_slave_spi_0 spi_0 (
		.clk           (clk_clk),                                             //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                 //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver5_irq),                            //              irq.irq
		.MISO          (spi_MISO),                                            //         external.export
		.MOSI          (spi_MOSI),                                            //                 .export
		.SCLK          (spi_SCLK),                                            //                 .export
		.SS_n          (spi_SS_n)                                             //                 .export
	);

	master_nios_multiple_slave_start_uP start_up (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_start_up_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_up_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_up_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_up_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_up_s1_readdata),   //                    .readdata
		.in_port    (start_up_0_export),                        // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                  //                 irq.irq
	);

	master_nios_multiple_slave_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	master_nios_multiple_slave_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                  // external_connection.export
		.txd           (uart_txd),                                  //                    .export
		.irq           (irq_mapper_receiver4_irq)                   //                 irq.irq
	);

	master_nios_multiple_slave_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                          //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.aip_0_avalon_slave_0_address                   (mm_interconnect_0_aip_0_avalon_slave_0_address),              //                     aip_0_avalon_slave_0.address
		.aip_0_avalon_slave_0_write                     (mm_interconnect_0_aip_0_avalon_slave_0_write),                //                                         .write
		.aip_0_avalon_slave_0_read                      (mm_interconnect_0_aip_0_avalon_slave_0_read),                 //                                         .read
		.aip_0_avalon_slave_0_readdata                  (mm_interconnect_0_aip_0_avalon_slave_0_readdata),             //                                         .readdata
		.aip_0_avalon_slave_0_writedata                 (mm_interconnect_0_aip_0_avalon_slave_0_writedata),            //                                         .writedata
		.aip_0_avalon_slave_0_chipselect                (mm_interconnect_0_aip_0_avalon_slave_0_chipselect),           //                                         .chipselect
		.aip_1_avalon_slave_0_address                   (mm_interconnect_0_aip_1_avalon_slave_0_address),              //                     aip_1_avalon_slave_0.address
		.aip_1_avalon_slave_0_write                     (mm_interconnect_0_aip_1_avalon_slave_0_write),                //                                         .write
		.aip_1_avalon_slave_0_read                      (mm_interconnect_0_aip_1_avalon_slave_0_read),                 //                                         .read
		.aip_1_avalon_slave_0_readdata                  (mm_interconnect_0_aip_1_avalon_slave_0_readdata),             //                                         .readdata
		.aip_1_avalon_slave_0_writedata                 (mm_interconnect_0_aip_1_avalon_slave_0_writedata),            //                                         .writedata
		.aip_1_avalon_slave_0_chipselect                (mm_interconnect_0_aip_1_avalon_slave_0_chipselect),           //                                         .chipselect
		.aip_2_avalon_slave_0_address                   (mm_interconnect_0_aip_2_avalon_slave_0_address),              //                     aip_2_avalon_slave_0.address
		.aip_2_avalon_slave_0_write                     (mm_interconnect_0_aip_2_avalon_slave_0_write),                //                                         .write
		.aip_2_avalon_slave_0_read                      (mm_interconnect_0_aip_2_avalon_slave_0_read),                 //                                         .read
		.aip_2_avalon_slave_0_readdata                  (mm_interconnect_0_aip_2_avalon_slave_0_readdata),             //                                         .readdata
		.aip_2_avalon_slave_0_writedata                 (mm_interconnect_0_aip_2_avalon_slave_0_writedata),            //                                         .writedata
		.aip_2_avalon_slave_0_chipselect                (mm_interconnect_0_aip_2_avalon_slave_0_chipselect),           //                                         .chipselect
		.aip_uP_0_avalon_slave_0_address                (mm_interconnect_0_aip_up_0_avalon_slave_0_address),           //                  aip_uP_0_avalon_slave_0.address
		.aip_uP_0_avalon_slave_0_write                  (mm_interconnect_0_aip_up_0_avalon_slave_0_write),             //                                         .write
		.aip_uP_0_avalon_slave_0_read                   (mm_interconnect_0_aip_up_0_avalon_slave_0_read),              //                                         .read
		.aip_uP_0_avalon_slave_0_readdata               (mm_interconnect_0_aip_up_0_avalon_slave_0_readdata),          //                                         .readdata
		.aip_uP_0_avalon_slave_0_writedata              (mm_interconnect_0_aip_up_0_avalon_slave_0_writedata),         //                                         .writedata
		.aip_uP_0_avalon_slave_0_chipselect             (mm_interconnect_0_aip_up_0_avalon_slave_0_chipselect),        //                                         .chipselect
		.int_IP_s0_s1_address                           (mm_interconnect_0_int_ip_s0_s1_address),                      //                             int_IP_s0_s1.address
		.int_IP_s0_s1_write                             (mm_interconnect_0_int_ip_s0_s1_write),                        //                                         .write
		.int_IP_s0_s1_readdata                          (mm_interconnect_0_int_ip_s0_s1_readdata),                     //                                         .readdata
		.int_IP_s0_s1_writedata                         (mm_interconnect_0_int_ip_s0_s1_writedata),                    //                                         .writedata
		.int_IP_s0_s1_chipselect                        (mm_interconnect_0_int_ip_s0_s1_chipselect),                   //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.leds_s1_address                                (mm_interconnect_0_leds_s1_address),                           //                                  leds_s1.address
		.leds_s1_write                                  (mm_interconnect_0_leds_s1_write),                             //                                         .write
		.leds_s1_readdata                               (mm_interconnect_0_leds_s1_readdata),                          //                                         .readdata
		.leds_s1_writedata                              (mm_interconnect_0_leds_s1_writedata),                         //                                         .writedata
		.leds_s1_chipselect                             (mm_interconnect_0_leds_s1_chipselect),                        //                                         .chipselect
		.mem_data_s1_address                            (mm_interconnect_0_mem_data_s1_address),                       //                              mem_data_s1.address
		.mem_data_s1_write                              (mm_interconnect_0_mem_data_s1_write),                         //                                         .write
		.mem_data_s1_readdata                           (mm_interconnect_0_mem_data_s1_readdata),                      //                                         .readdata
		.mem_data_s1_writedata                          (mm_interconnect_0_mem_data_s1_writedata),                     //                                         .writedata
		.mem_data_s1_byteenable                         (mm_interconnect_0_mem_data_s1_byteenable),                    //                                         .byteenable
		.mem_data_s1_chipselect                         (mm_interconnect_0_mem_data_s1_chipselect),                    //                                         .chipselect
		.mem_data_s1_clken                              (mm_interconnect_0_mem_data_s1_clken),                         //                                         .clken
		.mem_program_s1_address                         (mm_interconnect_0_mem_program_s1_address),                    //                           mem_program_s1.address
		.mem_program_s1_write                           (mm_interconnect_0_mem_program_s1_write),                      //                                         .write
		.mem_program_s1_readdata                        (mm_interconnect_0_mem_program_s1_readdata),                   //                                         .readdata
		.mem_program_s1_writedata                       (mm_interconnect_0_mem_program_s1_writedata),                  //                                         .writedata
		.mem_program_s1_byteenable                      (mm_interconnect_0_mem_program_s1_byteenable),                 //                                         .byteenable
		.mem_program_s1_chipselect                      (mm_interconnect_0_mem_program_s1_chipselect),                 //                                         .chipselect
		.mem_program_s1_clken                           (mm_interconnect_0_mem_program_s1_clken),                      //                                         .clken
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.spi_0_spi_control_port_address                 (mm_interconnect_0_spi_0_spi_control_port_address),            //                   spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                   (mm_interconnect_0_spi_0_spi_control_port_write),              //                                         .write
		.spi_0_spi_control_port_read                    (mm_interconnect_0_spi_0_spi_control_port_read),               //                                         .read
		.spi_0_spi_control_port_readdata                (mm_interconnect_0_spi_0_spi_control_port_readdata),           //                                         .readdata
		.spi_0_spi_control_port_writedata               (mm_interconnect_0_spi_0_spi_control_port_writedata),          //                                         .writedata
		.spi_0_spi_control_port_chipselect              (mm_interconnect_0_spi_0_spi_control_port_chipselect),         //                                         .chipselect
		.start_uP_s1_address                            (mm_interconnect_0_start_up_s1_address),                       //                              start_uP_s1.address
		.start_uP_s1_write                              (mm_interconnect_0_start_up_s1_write),                         //                                         .write
		.start_uP_s1_readdata                           (mm_interconnect_0_start_up_s1_readdata),                      //                                         .readdata
		.start_uP_s1_writedata                          (mm_interconnect_0_start_up_s1_writedata),                     //                                         .writedata
		.start_uP_s1_chipselect                         (mm_interconnect_0_start_up_s1_chipselect),                    //                                         .chipselect
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                        //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                          //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                       //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                      //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect),                     //                                         .chipselect
		.uart_0_s1_address                              (mm_interconnect_0_uart_0_s1_address),                         //                                uart_0_s1.address
		.uart_0_s1_write                                (mm_interconnect_0_uart_0_s1_write),                           //                                         .write
		.uart_0_s1_read                                 (mm_interconnect_0_uart_0_s1_read),                            //                                         .read
		.uart_0_s1_readdata                             (mm_interconnect_0_uart_0_s1_readdata),                        //                                         .readdata
		.uart_0_s1_writedata                            (mm_interconnect_0_uart_0_s1_writedata),                       //                                         .writedata
		.uart_0_s1_begintransfer                        (mm_interconnect_0_uart_0_s1_begintransfer),                   //                                         .begintransfer
		.uart_0_s1_chipselect                           (mm_interconnect_0_uart_0_s1_chipselect)                       //                                         .chipselect
	);

	master_nios_multiple_slave_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
